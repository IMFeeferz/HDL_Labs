module two_write_ports( input logic [2:0] write_addr_1, write_addr_2,
			input logic [3:0] write_data_1, write_data_2,
			input logic en_1, en_2,
			output logic [3:0] d[7:0],
			output logic w_en[7:0]);

endmodule			
