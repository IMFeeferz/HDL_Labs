module swap(	input logic [3:0] x_data, y_data,
		output logic [3:0] x_swap, y_swap);
	logic [3:0] XOR_1, XOR_2, XOR_3;
	
	assign XOR_1 = 
endmodule 
